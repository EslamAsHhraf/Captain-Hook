PK   {w�T6e� �P  o$    cirkitFile.json�ݎ$��&�*���d������
3-Lz/����J�-U����j��w_cDFfF�3�<�X��=huU��ύF���H����������<=�������׻O�����=��>��������Ǘ��?>w?���������_�T�<uc���<Z�|�{���N�yU�}��0�`�����������oG 6�~6.�~4l\�h���ѱ9p��gs�"�����EЏ�́���A?f6.�(��dC Sɷ��7�ld�7�ld�7�ld�7�ld�7�ld�7�ld�7�ld�7�l������,����,M��4|�Ɇ@|�Ɇ@|�Ɇ@|�Ɇ@|�Ɇ@|�Ɇ@|�Ɇ���o;�Ȃo;�Ȃo;��B L��N˷�ld���ld���ld���ld���ld���l������,����,����,����,��|������,����,����,����,����=�v�!��v�!��v�!��v�!��v�!����vz��dC ��dC ��dC ��dC�����ld���ld�������2=����r����O_���/Ň�!�;���矟�N__Aw�svV6N��Y�i���}�aHSo�G{'����G�bK���?�''�dw�g��@��~4��3$���ι��8�rQG�L�*��u֓N�c��0X~ONVV�VVeEف,;zde�de'�d١�C��(��3'7/+�Ň��I�=Ȫl���(;�e���좬�Dف,;��(ý�ݤ=xi
�AԪ�[S�oim��IV���{�U�Lq�H��u�D?��t�EÔs<�H@8���W*F��'II�R±,b���:L!c�U�SV.�w��8+7v�{7�1��-��+��irx"��`��ܕ\�+�i��iLQ	�c ���a~�[X~��eMuǮ��yj6���GT]�u)�^���6��4X�4����2�d��0�R>/,?��L��+������d��0��eAX~�	�a~e��p�_8`�����6a�	L��@�_��",?�G��+[s��'��$����ME��]d��0��JX~B��@�_��%,?��C��+[Є�'��a~e����Y~ ̯l���p�!������e0��,?�W�Z
�O8������&Qa�	���@�_��*,?�:6�B6���
�V8�����ʖba�	���@�_�-,?��C��+۸��'��a~e�����Y~ ̯l���p�!����M���s�;6E뇹Wc,f����L��Лa��Q3��e?V>�)*���	�.��@�_9��RkF���,6s�a�����Dd/�8�G��+gjPt�d&���һ���GLN8br��,?�W�@��p�$�����[��'1��a~��a�	GL��@�_90GX~��,?�W�����^������!E�g�L��
�	�%ݩ��W�:� �irܽ\�TDD/1��+'3	��p�#����3���'���a~�4,a�	�.��@�_9�KX~�'HA �x����.��@�_9;MX~¡�,?�WN}��p�"�������'���a~�=�����̓V���r�����JC����7X�v��pԳ�49<�/���E��+#RT�{�b?v*E�A�T�f�`�)�zH�rw��S�p�s��Ε�˃5�.���<�r��������Q��+��^m���ww>~yl���/ϻ��x��Vҹ�`8rˬW[Ϋ��}j�)g������t��ն�P�����3��2��E<{uYt��R��7�6�i�f���{��۱�]3�w{ֻk�L���TM�ݼ�v�w��۳�����Y�a�wd����5�F{7��kv��nVۚ]#�(������յގ�O���y@�e�:���z�&�1�<�>�$�Io�}3�́��!��Ys�\5�$����H{��D�1�\�g��o������w9����,�iTy���m��Y�]�gқ��h��3���<0z�6Έ��fV�����//�����M5{�j=��=_υQ�&F���M
T�����zw�Ŧ:l�w�F)�a㼻��Y㜣ʃ�����7�הJ>q��F4��7W6��B���f��8s�uM^Das|�u���0"75�ޢg=f�;kUL&�4�f�u�i�)��G5�!+g��uPS��΃��^We��q'뚬I�k����ɚ����Ӕ��v&G���a%�8ۚ�#���W�l\�┧>���~�?%RM�y��㎔���7��5����ZO��\�hқkM˩��\�V9��%����ͤf���c3���dm��ʛ��ʛk�Lz3+�\�gқy9�ʛ���f��`����ā�xs���4�qFO�,e�����pv���L�!(����ff��Ѓ���q`�|m��ƛY=_O>��'H�ד��ZO>О�'�+����� ��"�yw-���r ���L>�˕�q.�P�y�7W<��xsm��Rƛk�ǋ�3>�JF���2z��Q����7�z�JF�����:��+u�P��Q'=%�N,;�X���e�Y��9�Պ�e'�w��Zڻ��ђ�,3�xs��3�L��l섭�A�f���S:�ݘ�1]W�B�%ƛ�K��H{��D�q�S뚼����묵�k'���%��M��4v�=���\�/R�3��5y�إ���A�8 qL��^�l���L�]����ݜp�62���:j��ʢ�-2Ch�R���~rsu͇�&��S�~�POHLj/I�X=�2�/��#�`����T����Әz��P���qGz3k�פO���f��8Fn�頌W��dM�(���va����C���d�sʦl+	#�<�g#�v!Λ���U�H{�2*h�o��GZW1�\�WHz�;��R&$&�-��� ���'���Ќ�x=Bz��!=^σ������|=B�b��(k�}�Kƫk�}ګ��F��L�������"'�c����f��WSv�BgT����N�k0ֿ9�v�,$�G_h�{�k}���Ű6�T�1Ho�}3iGl5SH��z%IJ�ˉ�yFʫ�,�q�,�2���\Y��<���T8@Rź6�vs��6�����_ƛ���)zHbR��~�󠍚����	��vj|L�v�w���|3W�E��f�!�J,M�|�k��s�On0gi3�\���O?<����8<}yz����w��y����{�a�ݧ����}������#! ]�#! ]�#! ]�#! ]�#! ]22���tI.�0�%_!�HH��#! }Ȫ�H9�-g���6�n)$}H	q�� f����!%�I�~���B҇���8��p3�RH�pt�'1;n���>�%�I���s�����RH�pd�'1;n���>�%�I̎1;.��G�	q��F̎K!��bBḘ�bv\
	9��q)$�$�J��V̎K!!'1;.�Tn��$fǭ��B*7��q��V̎K!��DĒ�bv܉�q)�r��'1;���R9F���wbv\
�ܓ+�I̎;1;.�T�s�$fǝ��B*���-���q/fǥ��%�b�����RH�2F1Nr��r˛bv܋�q)�r�'1;���R�0N���bv\
��N&�I̎1;^CboA���F�p�W�=V��% �\����NU�+4�
M������}u2�ڂ+�r�K���nqTA}m��pŸ��\/o���@�Є�b7�мuy۷��\�Q�zy��8��\[p�&\����⨂rm��p]�������H`�UUP������
�Y-��*W�Es+�	���-��md�(�jv���.7�
Zh��[iXIٶ	�.wY�&la����`�&k�ڰ=�]^R�k���޶	�V�
�M m"�&l�۲��l�DcM�B�eOIٶ�Ț��6l�ޘ6�m�@�Іm���fa�M\ք-�a[�*��m���	[hö�j#�6qY�Іm�;�F�mVŚ��6l��6�m�5amؖ�|md�fu�	[hö�Il#�6qY�Іm�[�F�m�&l�۲G��l��eM�B�e�kٶ�˚��6l˞�6�Im�&l�۲���l��eM�B�euٶ�˚��6l�^�6�mT�ب\�M\f��e�M\ք-�a[�淑m���	[hö�1�F�m�&l��rVBٶ�˚��6l˙md�&.k�ڰ-gW��m���	[hö���D���α&la�����e�M\ք-�a[�DiR����e+l�a%e�&.sm�&l��rFM�m����V�6q�k��6qY�Іm93��l��eM�B���6�m�5amؖ3��ȶM\ք-�a[΢j#�6qY�Іm9S��l}���&l��r6X̷��V�J�Jʶ�z�o�5amؖ���ȶM\ք-�a[Μk#�6qY�Іm9;��l���蘏6q�o��6qY�Іm9˰�l��eM�B��L�6�m�5amؖ�%�ȶM\ք-�a[��l;�6q�
[iXIٶY/m�&l��rfi�m��������y}�۽ڋ�TN�݉R9�{'�[_�߉R9+{'J�t�(��w�N�������r<����uB�{��<i�8�t���s��������T���#���L���uÿ��>��90��Sc���8Nf9~�?�G�-�a��}�oF8hq�����2��A�C�L80��8�����8è���E���*�n��1u�=p0i����;C�K٨Ι�����aL�/�^͕����9/�P̖='����]e Ё	qVa�g]ҝ�9x���	&��r�	D��N�~���b�f��dIB�[ZGB	[ZGB���H(��Bv�Tn�ثu��f3V������c���ۚh0~k.��lz{9�a�sTyp����7�ה\��^C�kC��[f��@�]*t=(��Q�9�
G�0h���z�	e��0��V�����1��Y�"�YN�lf�os!��rIs��M��a���G��cv*;۫��>���N�z�LB�M�RP̖BB�[H�┧>���Y9?��5C�	>O��Q.1���E$��\b��(�Hj�	� ��c�S�R�A�0�t��U?�I�Nk��f��]WR((G�,�nJ��Ov�5�����k��u��)�>��'����Ѧ��!YNr��	�����:��]�Mǌ��阑P��h$����HB�t�H(��	e�1�iݦcF��t�h0f+�C��[���J��`�Vr���]?�<h�i��y7������g?�����5�IB�-�IB1[n	e;���lG��5E�P��IBَ")(�Q$e;�$i�vI�َ"I0��V�f����m��lf[i0�k9�4���9��jKFq�AM!;f{B�FBٌ�&�s6v� #P�0����)�nLƘ��m.$����4�q�0�ft^]�Ѝ�/r���L�6�&���ɪyrI9��>�i��k�\�%I(.	��j\��{����eZ2
�"�P�0�	Cx�� NB�L�P̖\H(�S5F'��ī���ⷴ��cߏaT��)��@��Әz����z��[_db��0�=�e�:|�����8��1׸�P���0ۀ�q�P�T���0Ø�:O'ݝ�ⳒP^�0����s�����+7O���8+c�hÀ_k�SD�D��/"�l��P6�D�fa		esY���9ÒP6�Dʦ�HB�tiZ�=	�`6�D�1��RsC��[�S4��(�#��'1�`K�*��e1��RkU����㔠�ʦ:� ���C�:�����A�4NL�˕Eʫ϶��Pl~���_p��r�	j��!�n�c�v�H(���LA�4�$�Mg����SP6��.w����	�k�1ŀ-��epX�o�	�V�H(fK�H(�}DB9.�"��(�}�F;v���ch2ͽ�1 *����朦�1MB��/���cXmԜ�\7N�u�S3������.ms!�|�������㷗�e����w��y����{�5م��闗���G~{�@
�hKE	��8a$�cV���>�FB@�`KD	�C  �HH�	FB@���0҇ G���>L2&R�j˙m1�b�[
I�BNb�Č��>F�2���7�p)$}ܤ!�Ĭ���B���#2�����RH���E����-瀋�q#fǥ��q��'1;n���>�,��$fǍ��B��=O2�����RH��K&��V̎K!�{��8�eR�R)bv܊�q)�rߌ'1;n��R��D����bv\
�ܧ!�I̎;1;.�T�o�$fǝ��B*��q�ˉ�%�����RH�\w1Nbv܉�q)�r��'1;���R9�Zl�G̎{1;.�T�I�$fǽ��B*��q�[ݔ[���^̎K!��S�8��q/fǥ��y�b���x��RH�|H1Nbv<������g�J��d@�&\�	W��8GTUP�-�B��qq��4��\[p�&\���^iTA���
M�b��D��+D$Ђ+4�~P�.�s�@�Є+�(M亸�AD-�B��qq��4��\[p�&\���iTA���
M�����Ҩ�rm��p-5�m�6W�Іm�mn#�FQW���M�m/hy5amؖZ�6�m}5amؖ��6�m�5amؖ��6�m�5amؖ=md�&k�ڰ-{1�ȶM4ք-�a[����m���	[hö�i#�6QY�Іm���fa�M\ք-�a[�*��m���	[hö�j#�F+b�����e�M\f��eM�B�e\ٶ�˚��6l�^�6�m�5amؖ=�md�&.k�ڰ-{+�ȶM\ք-�a[����m���	[hö�um#�6qY�Іmٳۦ0�M\ք-�a[���m���	[hö�n#�6qY�Іm��F����+���l��̶�˚��6l���6�m�5amؖ3�ȶM\ք-�a[�Jh#�6qY�Іm9�l��eM�B���6�m�5amؖ38��ֵ�˚��6l�Y"md�&.k�ڰ-g���m���	[hö���F�m�&l��rFM�6�I�h+Y��̵��\���	[hö��F�m�&l��r�Qٶ�˚��6l�Nmd�&.k�ڰ-gQ��m���	[hö���D��M\ք-�a[�k#�6qY�Іm9㬍l��eM�B�嬶6�m�5amؖ3��ȶM\ք-�a[��k#�F�|4:�M\���e�M\ք-�a[�2l#�6qY�Іm9���l��eM�B��l�6�m�5amؖ32��6��˚��6l�Y�md�&.k�ڰ-g���m���	[��}�*z��~���f��.���zTnt]�r�j�0�D��M��r��N��9�;Q*'o�D�����r��N��y�;Q*'H�D����W넔WF{k�����ժ{ad4�v��^�]�FF�k�q���2Z\��r/�����#�ŵ���hq�^ý����n|���O����!ʥlT�LP^O��0&��m���"�es@�P6�� �g&|�%ݩ��W�:� �ir��\H(�r!�lʅ�"#�M3CBٴ2$�M#CBٴ1$�MCBٴ04�R^����h02�����`d4x���Y㜣ʃ�p.@�d����䢎GMI(��mu�|��
]��iTy���m��Yos!�lr�۪��V�8f�;kUL&�4�f�#NBٖK��s��>�|�S��^��y��0�D�E���$�l���)O}R}�r~�?%tk��E|���m��P6�BBٔ	eۡ���aD�&ӫ~6���֦�	�@�	e;ԡ�lG:�M�x]��N���e�<�����6�^�ڰ-ʦ\H(�r!���es^#�lNk$��Y���阑P63ʦcF�:!���mǌ#��ێFF�����'��:�14��"�U��g���zBIA���)(�n8e���l;��m��"���Q$e;���lG�$�R^�%D�$�%D�$&�����~�-�Q5��<�i�	�	e��'�s6v� #P�0����)�nLƘ�#x�$���4�q�0�ft^]�Ѝ�/r���L))R
�&���ɪyrI9��>�i�_wS�	r!�lG����OjP�%C��+�
���0�w�蚂"�e�:�P6�	e�6�P6MCǾè ��SR�3�Z7�1�6ρ��$��>2�KS����2�Y>��z`s)��6fp4NJ7�J�XaSA�������8�����q���Ӭ�4���>�0�ך�0�((2\��e{QP��es�P6gXʦ�HB�tI(�N"M넔WF{��D���n;�4&8�Q똜U�b~ѥ
֪��1���)��$RP�3��-@���н�Ψ�q:v�;��H�BBَO�Pl~���_p��r�	j��!�n�#!-IB��*QP�#%
�v�DA�]�&��+HN�1b�[S�ఖ���P6�����G$��>"�l�	e���h��BR1zM��W�ևX	�NksNǌ��l�S�a�Qs��q�8���N�ަN;�;	�#����������������>����|~��=��������ǧ�qz������\�Y�?���f`�sp�lYu:�7ƛu��ĥi�r��ħ9���7��]چ%�ʨ"�hp�]y3� �#m�%��7S�-YEG�wSg����Zoj�,�����ȫc�;4�5b1�zE�%漺2eR�k�-p
�8o�X4��`�&��6���+�5iӊ~8�ޜ7�L8mݞ�f�����V��YgYP������-4��eֻo5��n�[{�yHD����k��f}7��Y�V�9���Sl�ys���Ţ�7W�8�����'_V�L,���8Բ(��9���o��3�8������Dz�Tֻ+.����}7s��t7w��/fV�"{� .�Qâry^	G,L���y]�D�fv���L*N���
b�%�˳d9�>w�h�q�!�IzJ���T+V�L���T�U�L���T"r�\K��1|3�ζ�fZ�"���暴iՌ�D%�����t⽚�ϬW3�m�%VnJ1�b�6�S��`��8�̔����*���P����<χ�m�Ԩ��Q~�c��yk�MZ�b�Ϥ�;KRb�!�
-J$�q
�j.�p�S�����b�ZB�V�)�l���B�ʛ��[_�hb�*k�e҈'V���\��O������O�6����q��������y�T^�"����`}�	0k?��%�W	|�JЫ�GA(��u��.`���Y%z���)�J��Ԍ(������j�Q����5/~�:Z
�rZ
ܪ���{��pkl�C��l�w��,�w(6�`�7�����|$j��.���|�zd>fY2� �:Y`B�)P��*P��,P�V._w׿K�_������NT'��nE(p�###N�����[���M��]�V�_��=
�����|̲w>f��Uߣ�zV�;���%�,��K�Y�7E�y
�:���H�
��`��U���p_��~_�#����R�!��|!I���ҵ�|F�%�\3�	��������Ko=�kʏ��#�'�*��5�*��C�*��Q�O��_����&���'���(�/�|���[*��wV�		o��N�;�hf)��-��u�'��|�g ���v}�j��#[n�w،��PP��DH̭)�Ñ�C��Hz��UF�c�����;l[iF��{�z��;lbi�Խ,W	|�--|�;[���7��-.�����O��^������ߟ����Ǘ��_>�w������y���	ے�^�~�H/�!��D0Y�!��� &6�>�;�d��Ї{�,��p��B.(b�`C��GLl}� �ɂ�,1Y�!��&�ْ���S�~���c��S\6�(Co����� `H�e�H���-c��Х��C��{��Х��C��pH���|]*X�<���|]� �y�S#`O�������F���1t�d�%���|�!`O��C"���V���1���=�c {��@����<�)y�S>F)�H�	�S'`O���X���=u���Q�gx�S'`O��C���1���=�c {��@������=�c��j���S>���|�!`O��CbJ��z{��@����<�)y�S>Fْ!�P)`O��=�c�-h<���Ow��?'[H��g����=K��˔.��;����@��Y����̆:���@�.,�2?�
��
��,?��������d��0������c����\Е�gV� ,?Y~ �O?Fa�Ea���a~��������8t��Dę��1_wv<�ّ�K�\_Y688���a��zSZ���x#�\�Z�C�A- %�
aA@�J2�;��ifJ@:�Y�J@:���F�!H3<?REF����\--3}&LVs% �t�#���?$#C�@G�!H3,���2��n��4�R�/-Cِ��4òA:#.�3i�e����a� Ͱl����t#����+�2�^�f�˶iJ�-�A�a�2$-C�a� Ͱlw���t�"����Z�2��S��4ò�LZ��q�0C�fX��I�P:Nf���>�R�8E�!H3,[�e(�3i�e[����a� Ͱl	���xݘx�t�b��+�3i�e+����a� Ͱl#���t�"���-��2��S��4ò}[Z��q�0C�fX��K�P:Nf��o9�)����bYj@�0��J@:lq�a�0C�f��2m�EF_F��Q�0�r��ZJG1�A�����Z2�v�b�w�H5N:�q�A�0C�fX�򐖡tP#���sH�e(�3i��iJ5�A�a9�EZ��A�0C�fXή���^|f����^�:�{U�tP�$,(#R�/�3i���#iJG1�A�a9�IZ��a�0C�fX�������}����a��[�t�"���㾤e(�3i��2iJ�-�A�a9fMZ��a�0C�fX����r�n� �,	ʈTz-&H�-�A�a9��Z�EA:�Y\a����!�{��d>�84q���cw>��&��Ip��[w>�8su��Rw>��p�[\��v�7I���
KB��gx�q��_��-�4��U��-l{��z�^������:n2� ���Vnr��-U�r��Y�<p�g�*,�--�a��/�X���5�{��C��c9>t��-Ǉ�\���_�P�ߘ����(�\�Fu����Mc�y\�ӵ��)pKv��n9xu��!�-Ǯ���:0!�*L��T���l�N�4�~Mvv$��qحȮ2ד�Vd�pWfz��K3W�[܊���-	�_Kz~qv���g��U�+�+�J�EXQ�ʼC�[��ʼC�[�۵y����Еy��wő�Y㜣ʃ�p�A�d����䢎4���x'����5�:M��A����4�<�YMZ:��f��	��|F|H�����1��Y�b2!�y6�_��21��V����`S�~�{5�]������j0��Co�)�v��������b�Ip+�zŰ�.Ny��;���#�)�76�.������TdG�[��TdG�[��T�������\�V9������ͤf���1��d5Ϛ�2*j�?nE�*]A�[ѻ��x]��N�:���<����Ȏ6�^�ڰ�w��%���]�gIp+zW�Y܊�Uz�w��$=�Qs�r�j��<	Iz���Iz���IS�+�&���IXQߊkH�[�ߊ�J�[I�W�D�R�k)6�Ws����A�N�Q�n�9:Q���~���_�j�%neb�������S�V&�ZҀw-��<�ԅڤL�[�ڤL��GS��GS��G�T�ZM�G� ��o=�Mã�ix��7�ڂPN!>�a�Dے�uPS��΃��~-R��w=�����	cI�]��C�t�1c�n5���W܊_Y�&q��8cDn3z�.�S�S�Ǻ~tsJ&�k��;��v�`�d�<�����鳚�_��)�k����8�2P#���I�v@I�(���B���'�&w�R��<}��4C5a��V�+.	n�ê(	ni�\��cߏaT��)��@��Әz��6j�A�[Q�
;�4���.�-Ҙ���m�� 6�q5�UcG���΅�󓇀]@%k,�0�)���Ʈ2]��VFEe����Y�8y��iV}gelmP�[aǂ[�]�cIpW��Hϯ�ZV�����U��])!=�1 =ŷ%=ŷ%=ŷ�)۵�pŷ�,'�Z�oEa+��JpF���U�5j��ʢ�[�1:t�Z�r?�~�8g�y��i�G�q�A��WSv�nBgT�P;ȝƹl\c�k��%;_ͧP&�g�	?6���s�؍C���p�#=�2��"7
�kNz~ep�?
ܵ������+Sg��	�+HN�1�[S�����Y��Wt�2ב�V
5+�H�[�����$��L�+v��ҕ#�F;v���c 5ͽ�QK��ή�9�5��fHp+=[�X�O}�Qs��q�8���N�ԧ#�ޭ���ؑ�V��������������>��Rdv���we,^�S��e.*S:������X�=,�����!�zH�r���!�t��;���a�鰎uXP9,�"�C����l�����Մ2�%}|�R4!���NJa��;*�]�p� �|���5�U�Q�W����>HY{��1JJP�����YR2qgP�cgP�U�zHȊ�� ����)������7lq] 8��]K�k���VW{�2�_�L���H�?<���/�9���R��G���\�W����Sjz������2�C�W �$c9dx��K2�B�Xcȩ���C�ʇx·T��XUz��0wp_�q��J�H��q�U���Yt���K:�E�UmW�dVi�ʈ��tB�y]O�7-���b�,�͊�ڄB,~�,�s�~�R���Eᜢ!N�l^�S��JmV$��r
��dj3��SĶ$S�Ph�Ҝ��%��tB+��Ԅ-Ș����qe-eÛ�8j�:���6֐Z�jMmn�npfU�-�Ԧ�N���LmJ ����X��Yb��N���L�7�p
�dj��X7Ʃ��l�X~H͊7Vpj�8U�<�l� �e0k���b��3�����iy�-kk��a�5�M=_��K�w�,�U�<���<vg�-�U37���<vnk���Z]:u�RX�əx�KX෺�fʉe��PN���Cj�N,{攞r�j9eLK!Ԧ b�*��sA��& b�+��uI�6�Pk�n�F�6�d�B�v6y�M5�D+�eY�����fBb��թ��&B��9�%�Z�A�yq����5�M4Ľ�U�-w�%��q���r��,���}8��k}^�����<��n�_�����<v[��MX��>N�"�z�!���XYȩ���.?�Z@+����.�ԦEb�0ø���̓ĺ`�P�[�f܉e�,r���z�����K�O_Jy��������^�S����O��ɼ�d�?�ן��'���[��_�˟��Oa�S|�).J�?��O�����	NҀ�8�MKy�I��K��I"�	�DK��I&�
��K���7��o8I�"���`)3s��Y�̼��R.�$���9��,�bNr1K���\�R.�$�"������������ٓ<�R����v����}v�}��}v��N}d�}d��R����v����iW0Or�K���\�R.�$���;��-��N�����ެ�Rf�$3���;�[�;�ŭ����]y�$3���;��-e�O2�K�����Rf�$3���?��/e�O2�K��7����?};���˗��y����{?���|��Rf;��,Ɛ�����t|T���/��r��n��6�~���.���O�{~�yz~�<v�������?�����Da|��\�^~������/�o�GL(�����H����OO���'��}��/�&��������}�Lo��<��_>?O�ݧ��s����^~y����������_�� �>�|~B9���{����,�~���;��i���ZE��i��Ko�_���0�?���}�ϐ6���==ƾ�L�?��O/��������ځ�W&>|��3A��.?������yCk�x���ix�����ߪ��6�{"�]�~oi5/����������]���Xi���
�7$,G��$�H�J��)XHXn9bVZ��xYiIX��u���V@²$,w������?�_�����ӿN�ߎ��A�̝���������Ͽ|~�O��:�R�����T69�6���2�!��ؔ-�T�9+=D�� �1f0����i���r;�"��z*g��-��5e���gS��u&��Qɪ�\z�?�����O���x���V����x�^��̢��p����� ��/�'�u.��Ѕ��]�R���y,JS��Ns��9�^���b�PrQ3����F����5&�׏�X��=�d0B>~T����]0)Ր g��C�t�z���.D8YE�H����r��_!e����Ѫ��{�WF�y�!�o��u��{��h r��,JFbr��ht���/t���7�������4p�r�ws|��$*�����Z3�hɇ�����
���G0�u���m@�ơ�q�-��T���8���~��glT�Q�8�s{�����O�MO�q�9�@��Hœ�1�p���4��˯����tCV)H'&����Ôp�S�&4
>���"��0���sx��?��0�.��7OHga�+�$�����&�#�p��[�"�������sU�:h�"�'T���ha@u��¯�*���w٣��p�I�}\�䗟�0%p���P����Y��9����;���oP��c���C�	���^c��HG������������b��E�+�W���O�p�FG�菙��7��tH����U��
�SV�-�'��*���B��|Q���U�|��_����ܹN}�D���#���t�ݹWo�~�}��?n�O:��QYC��O�a��?���4��=D�`�����n}��h�`�� �O#q�:���]�!�e�%1];�kqF�cB�]�=�����-W�N�A.�����zmf0�mfХ1%mqJ����bG����u<ܛP�	�+�_mf�L8�ϚW���g�	��J.�7�4�������������GoݵV��^�Z~ޯ���WC�|�'C�f��B��m��,��g{�lx����}�#�����4|4�?���xOS'8���|��èvo��-��N6_�_����X�ż��-��2���p��ׁ�j~J0�����(������A�0��~�:�S�4���'�:�O��E��_Cz~u�)���y�Jn��I�"R}���c ���́��jp�o��S(���|Gm�\u �yI�Q����Mʿ���h ���(,���e���2%N��A减�����x��[m�O*t6Ã�8w���N���'�㿠����!L�Ai�q0(�@f�a�}��L1\��t���Ƨ�|]HO�aQ�>ù4JX����o�a0 !'��q������>��'��e���ù���Y�`:����4�A�!��g~t�H%S��%�*(_��`�K6$���7S��A|Iû�vx=��ɫʕf�!��V�0�E}�����k�9:���Q�8s���[h��ud� F
�`O	��i�4Ƶ��S����P�nFp؜_t�gLs��4�|��Wal��zZ+�	Av��tn6UEt�Ȱ��-����f����;8T���Gk�w��+	��J6soP=�u�X+m�sY��Vi��i��0$��q�r�#��Ns�����+�?��t�����k�MBSJu�ǜ|�7Ɵ��5^��t>>aqY�{J����/N��1�ת�XRP�-�C���p�)<�`�CL�W����24�5>��9ax�̮�V�����Lzp(�|r��zz@�O�Ն��u�ѿ�~�.��^�S����"��^���!,��Ʌ;5�;�y��+�R�w�\(!������+͌�~��+�����G��Y�ᵙ?�� �o�k��>�򯝘|���G@[�=����x���/\��u�tq�'|0���16���Ȟ�H7c���p��V��o8`q a�w��_����b��hHE|��';|�B��Q��ٓw"Q���R8�s_�{�dF�f.H׻�$�{&r::�� ��1�'�}�1w�� 8��)���,~�h^ILOk�����8t��|,�+��8�+H��k�H]�]<�])����i�*an����!v�9V7��4{��	�,(���hp�|�(�Q��U�mNw�bW��v�x���tX:px�{*���B`��������k�utps��h��tHC8T���9��7�_~��>���U}H\} ]�EL�ۏ���љ> M�)
O�|z�򄂻S��⇔~>���:&����<����B��c�é�d��h�}9��������/7	����v���������/�7vӷr�����j����w��p��5~c�����K����_;~���+} ���W�hw�������$5�����������ﺗ?����?�ᮜ�������r��ʿ~�}���=��eh<�;;����Y����Z3�nkf�C����T���g��k��o��ҟ�������kd��N��F��Fa�Q�"����\����lyU�����Қ�+�����VU�=��JoF�n=��I�r���mE�D��}������:Cnfώ�xW�����ff���:4�N��:d�tH��!-�Cog=\�!Z��r\�+b3�a�<�L�!�E�$��;Jס�:���Nz��{�'V'�E3�>L������]}�����+϶��[-�񏥴�o���`�Qi�-�[3�/�#���A*gF�����f�����&����v뱰F����vj�ewV4r������ՏRڵ�?J9v��Nʱ>߹tS3c֛�5= �[U����s���բ��F��u�d_�NW�}*���2t���fO�v8��h�'}6wR���	�U�zr���TD�$�H�|0kx�u��o���C��ጲ��Nk��Ss���Ҫ��Q��z8A�H���d�#I���Iw��(�$o��f����Mmv~VlU��j�(��U6ZN�֙QZ��Y�=���v:}ќ����U\�xYҚ�_\S�e�ue]2aU6Z�֙;ַ��S��V���v�u-�6[7Yq�����Ue[��Y�n�ԥT�U���f��'�ܤT�ޔ�0gf�1�/۟���z��r�[�ZW���!ϒ�!8��= tnb�q�
��j�' �9�|h��78UUcѪf5Ҝ�S��Kj��p�Ξ,�j����N�x;����]��V� �e�<�+�U��ċ�Z������V�����RE�10{V)eUq��h���S����[�����a<��-�!�d%i1�O�P;��;�I�ϛ��	�3��J{�j��,��z�Z��)�1y�%�뎑����m�nBW��c�#�J�d�q�q}�Q�����T;��rPз.�2�R�Aktw*�� _��a��|R����Q�ڨV��M%5���΂�3�F1>tv������C/e[1>筌]+Ĺ0Q�V��p���f�]�ݙ˶��ǣ�?��\�Z���s�-y���D�ɕ�A;b�Ԥ���X9�s����y�J���j�ͥ�+Ǔ4wG����h��]͂G�YI'.�Sth���������>~<�����e8W�f�bڞ/�Rۡg���R��*+�!uS�T� �F;29;�I��M���C��jt�L\�ή̸�F�vk4�� ����ذ������M[V?�h~T��S�?�$%T�ָ�w5[74i�������o�.�O�֕��0S��h�)�V/��I�����]*����W���l�lyO��.��uhb��Q[Y��.ZU�OI�JJV4����M7E�+yv�D��Q���?{a%I��zhr���Vg��Ww�j]q�w���dݧ�V\�O'�����\�Hj�uSj�-.�Yp��e�ue��<��mԔ����I�Ň{r�;�4m��!I<�:�Y��\����c<�H��υ8��ne�--�@�h���Ӓ�/^J�J�sfj�I}hYI���p[wP����*x.�Y�5;S�Y����me*/Ռ�l-�x���f�I=��썒�����{Gq5)m�-�xv����}�l�y��L�ѝx��W�h��z�å	%63��m\4�hc�b��i�HR�HD�&������cE/[�&�s�Glf�sG�Go��Ҽ��E�Z�#z�ԝ��N��(WZ��#9ô��^��K'�z����R���9�%�h��K%���)�6jab�pG�l)!�~�]���R�-%��n�Q��NQ�B��ew�J��y�0�UUwլ��-�IR-io������g/?\?��7c>�a��Z���H��U���o􏩈7T#��'%4S��?�����E+b��.��1�E��=�<�2�"s�m�n��-�"N!���y�D�ւ�{���=�I঳S�9[$1yu�.��j��-�����W�;_�#�򔕽e�J�e2��b��ʞ��&��w�E;SZ�WW�.ԑڊr�6��_��r���V�:�e�Z�h3������f���j���3JkV��.Ց؊r���_�Ǘ�Hk�H�v�J�o�M�Q40q�&{�
F&k|���pѕf��/Ԃ�j=kmù�%���w�d�Z�,C�����>�E97t��=}_�?ҕuWI]]��;����ԝ���VP9�����V��WR�]�l��a�Fc����~��e���y~3�U���Ԉh�&f�B�
q�qN�rb��M�T^��q�����z�k�Krh��#��V I�����#�����j��NS���_�S������}㉉]�z�*����Y��O��z`s���q�>�2� .OI�΀�ܜ���<�]5;�l�v{{<���p�E\�M�hכA�M����ι����_��f�B��S����f�P��YO:M�ɸ�;	'�Щ�c���q����N�c����
 /�	Z����{�l�f�]�!4��$��V�H�xG6v5)sS.V��8γbc����)(����vD#�KA��k'���%��M��4v�4�Shg �A�:t[AvP�227*��5s����_]A����-�q^K�*;��D�qV]�V�܏�<��]g.�Z���Y�xS���&�]z�p�{�-�W��)3��T7G�svV6N��iV}B!�G�I�Q-��=Zm݊ *Ycq؇aLa��]�ѩQ,��^EBO;��d�1or�[��b�E�J�r~\0��"X+b����$� �ʐĿǇ�S�R�۬�e�����P�p]9*6�׉�|Ɨ&tUO/��Ւ�zjZ�6<�j;�j{�Ie�nJ�a���"G8\j��u)[��C/��_W���!W�f��.�1��@cl-�D�eR;���p�R����F�G��ו輙�D�p~��Y庖K%"^ײ+;K�(��쭫�;�
&g����G���S.�9���Ɩy�B�ΛU�*w��!6[dq��,\o%q<3��d��o=�w�6v���\K�x�T]�Λ��=��|�6[��}�a-J,H9YY3��0:UA[a�W�lH�H�ͮ>���c4�,*�.�$I͈f'O�#�ă�I�ҋ���w��v{�؟9is��i�*�o^�=��7�MJ��V�z�Ż�NJt����'�K���`�y��2��j���u���Hj���e�M偓:r��һ�D %ݻ'�H�&���-�X�:��6�7#�|p��Y�Cu^Am�+y ����vԄ�e#�+�r���Chɋ�������^z������fD�]6�e�'��;��)��m���p�Z��~D7�wS����\�=gjҹ�yL7�Z<�xDQ2�A�́��yQOJjU�1��]"ߘ�#�"�_6�{c����d�
����e
0&��Zq�l}��ˣ�H�*y"�[j���D�7Y�n�ճ�����7��v�1!��:vѬ�<��c�͈9 ?�Lum��σ6jƨS�n��Gl�����i�{w}��;T��YH*F���4����p�˓���Z��A�0w�`�ۏ>w T�v�t�7�[�W@A���Ք�tF%��ұ�����Q� �A��*���8���V��ڝ_,_Wj;�"�!�IZ��L�y�Ԥ��|~JX��,�U�99���\A��MڃW����!j�~��ԅ�Tem���wY���{)���x�.�Ҿv��鞪���F����*Ȏ4�jR
r[f1��2������z���3�=䷄�5���BI��d�eG���&�a����q%��b�o5��l�+[��ņob�����2�h%��!��l:&ߘ��AU0R^a�[�B��e�k�E;]���y�;�]�L�Od3-��D�����v��$�1�RW��v��&n/.�!��,l^�V2?�����|����u/����˷�OE����O����}�/O�����o�������_PK
   {w�T6e� �P  o$                  cirkitFile.jsonPK      =   �P    